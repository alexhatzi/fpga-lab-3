/media/alex/secondaryLinux/FPGALAB/lab3/lab-3.srcs/sources_1/new/ps2decoder.sv